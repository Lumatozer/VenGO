package print

struct Hi {
    a->*string
}

function print(a->int)->void {
}