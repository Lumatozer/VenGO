function mult_2(a->int)->int {}