package print

function print(a->int)->void {
    
}