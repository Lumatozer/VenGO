package time

function Time()->int {

}
function Since(a->int)->int {
    
}